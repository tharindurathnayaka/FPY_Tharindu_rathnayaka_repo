module jtag_tb()


jtag_intro jtag_intro1(CLK_50,RESET,LEDR,R_IN,M_IN,PC_IN,INC,CLK_IN,INS_IN,CLK_INC);



reg CLK_50,RESET;












endmodule;