// jtag_uart.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module jtag_uart (
		input  wire        jtag_uart_0_avalon_jtag_slave_chipselect,  // jtag_uart_0_avalon_jtag_slave.chipselect
		input  wire        jtag_uart_0_avalon_jtag_slave_address,     //                              .address
		input  wire        jtag_uart_0_avalon_jtag_slave_read_n,      //                              .read_n
		output wire [31:0] jtag_uart_0_avalon_jtag_slave_readdata,    //                              .readdata
		input  wire        jtag_uart_0_avalon_jtag_slave_write_n,     //                              .write_n
		input  wire [31:0] jtag_uart_0_avalon_jtag_slave_writedata,   //                              .writedata
		output wire        jtag_uart_0_avalon_jtag_slave_waitrequest, //                              .waitrequest
		input  wire        jtag_uart_0_clk_clk,                       //               jtag_uart_0_clk.clk
		input  wire        jtag_uart_0_reset_reset_n                  //             jtag_uart_0_reset.reset_n
	);

	jtag_uart_jtag_uart_0 jtag_uart_0 (
		.clk            (jtag_uart_0_clk_clk),                       //               clk.clk
		.rst_n          (jtag_uart_0_reset_reset_n),                 //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (jtag_uart_0_avalon_jtag_slave_read_n),      //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (jtag_uart_0_avalon_jtag_slave_write_n),     //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                           //               irq.irq
	);

endmodule


